`include "alu.v"
`include "datamemory.v"
`include "lshift2.v"
`include "fsm.v"
`include "mux.v"
`include "signextend.v"
`include "regfile.v"
`include "dff.v"
`include "instructionmemory.v"

module cpu(
  input clk,
  input

  );
